program test;      

 //LRM keywords $scope, $list yet to implement

  string s;
  initial begin
    //$scope(s);
    //$display(s);
    $list();
  end
endprogram
